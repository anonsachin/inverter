magic
tech sky130A
magscale 1 2
timestamp 1766844613
<< metal1 >>
rect 24722 4356 25122 4362
rect 25122 3956 27660 4356
rect 24722 3950 25122 3956
rect 26492 2906 26498 3086
rect 26678 2906 27268 3086
rect 29388 2906 30362 3086
rect 30542 2906 30548 3086
rect 24260 1510 24266 1938
rect 24694 1510 27358 1938
<< via1 >>
rect 24722 3956 25122 4356
rect 26498 2906 26678 3086
rect 30362 2906 30542 3086
rect 24266 1510 24694 1938
<< metal2 >>
rect 19031 4356 19421 4360
rect 23896 4356 30197 4471
rect 19026 4351 24722 4356
rect 19026 3961 19031 4351
rect 19421 3961 24722 4351
rect 19026 3956 24722 3961
rect 25122 4067 30197 4356
rect 25122 3956 25128 4067
rect 19031 3952 19421 3956
rect 26498 3086 26678 3092
rect 26498 2681 26678 2906
rect 30362 3086 30542 3092
rect 26494 2511 26503 2681
rect 26673 2511 26682 2681
rect 30362 2673 30542 2906
rect 26498 2506 26678 2511
rect 30358 2503 30367 2673
rect 30537 2503 30546 2673
rect 30362 2498 30542 2503
rect 10409 2352 10799 2354
rect 14857 2352 24638 2353
rect 10403 2345 24638 2352
rect 10403 1955 10409 2345
rect 10799 1955 24638 2345
rect 10403 1949 24638 1955
rect 10409 1946 10799 1949
rect 14857 1948 24638 1949
rect 24233 1944 24638 1948
rect 24233 1938 24694 1944
rect 24233 1510 24266 1938
rect 24233 1504 24694 1510
rect 24233 1478 24638 1504
<< via2 >>
rect 19031 3961 19421 4351
rect 26503 2511 26673 2681
rect 30367 2503 30537 2673
rect 10409 1955 10799 2345
<< metal3 >>
rect 201 4356 599 4361
rect 200 4355 19634 4356
rect 200 3957 201 4355
rect 599 4351 19634 4355
rect 599 3961 19031 4351
rect 19421 3961 19634 4351
rect 599 3957 19634 3961
rect 200 3956 19634 3957
rect 201 3951 599 3956
rect 26498 2681 26678 2686
rect 26498 2511 26503 2681
rect 26673 2511 26678 2681
rect 9845 2350 10243 2355
rect 9844 2349 10804 2350
rect 9844 1951 9845 2349
rect 10243 2345 10804 2349
rect 10243 1955 10409 2345
rect 10799 1955 10804 2345
rect 26498 2343 26678 2511
rect 30362 2673 30542 2678
rect 30362 2503 30367 2673
rect 30537 2503 30542 2673
rect 30362 2351 30542 2503
rect 26498 2165 26499 2343
rect 26677 2165 26678 2343
rect 30357 2173 30363 2351
rect 30541 2173 30547 2351
rect 30362 2172 30542 2173
rect 26498 2164 26678 2165
rect 26499 2159 26677 2164
rect 10243 1951 10804 1955
rect 9844 1950 10804 1951
rect 9845 1945 10243 1950
<< via3 >>
rect 201 3957 599 4355
rect 9845 1951 10243 2349
rect 26499 2165 26677 2343
rect 30363 2173 30541 2351
<< metal4 >>
rect 200 4355 600 44152
rect 200 3957 201 4355
rect 599 3957 600 4355
rect 200 1000 600 3957
rect 800 43526 1200 44152
rect 6134 43526 6194 45152
rect 6686 43526 6746 45152
rect 7238 43526 7298 45152
rect 7790 43526 7850 45152
rect 8342 43526 8402 45152
rect 8894 43526 8954 45152
rect 9446 43526 9506 45152
rect 9998 43526 10058 45152
rect 10550 43526 10610 45152
rect 11102 43526 11162 45152
rect 11654 43526 11714 45152
rect 12206 43526 12266 45152
rect 12758 43526 12818 45152
rect 13310 43526 13370 45152
rect 13862 43526 13922 45152
rect 14414 43526 14474 45152
rect 14966 43526 15026 45152
rect 15518 43526 15578 45152
rect 16070 43526 16130 45152
rect 16622 43526 16682 45152
rect 17174 43526 17234 45152
rect 17726 43526 17786 45152
rect 18278 43526 18338 45152
rect 18830 43526 18890 45152
rect 19382 44854 19442 45152
rect 19934 44854 19994 45152
rect 20486 44854 20546 45152
rect 21038 44854 21098 45152
rect 21590 44854 21650 45152
rect 22142 44854 22202 45152
rect 22694 44854 22754 45152
rect 23246 44854 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 800 43046 19218 43526
rect 800 2350 1200 43046
rect 30362 2351 30542 2352
rect 800 2349 10244 2350
rect 800 1951 9845 2349
rect 10243 1951 10244 2349
rect 800 1950 10244 1951
rect 26498 2343 26678 2344
rect 26498 2165 26499 2343
rect 26677 2165 26678 2343
rect 800 1000 1200 1950
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 2165
rect 30362 2173 30363 2351
rect 30541 2173 30542 2351
rect 30362 0 30542 2173
use Inverter  Inverter_0
timestamp 1766062202
transform 1 0 27626 0 1 3512
box -700 -2000 2056 800
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
flabel metal4 800 43046 23716 43526 0 FreeSans 1600 0 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
